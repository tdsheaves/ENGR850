module arrays();
int l_h [3]; 
int arr2 [8][4];
l_h = '{2,5,3,6};
initial begin
bit [31:0] us[5], dub[5];
for (int i=0;i<$size(us);i++)
us[i]=I;
foreach(dub[j])
dub[j]=us[j]*3;
end

 